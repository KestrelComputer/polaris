`ifndef POLARIS_ALU_VH
`define POLARIS_ALU_VH

`define ALU_ADD		0
`define ALU_SUB		1
`define ALU_SLT		2
`define ALU_SLTU	3
`define ALU_XOR		4
`define ALU_OR		5
`define ALU_AND		6
`define ALU_SLL		7
`define ALU_SRL		8
`define ALU_SRA		9

`endif

