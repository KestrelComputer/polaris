`ifndef POLARIS_OPCODES_VH
`define POLARIS_OPCODES_VH

`define OPC_LUI		7'b0110111
`define OPC_AUIPC	7'b0010111
`define OPC_JAL		7'b1101111
`define OPC_JALR	7'b1100111
`define OPC_Lx		7'b0000011
`define OPC_aluI	7'b0010011
`define OPC_CSRRx	7'b1110011
`define OPC_FENCE	7'b0001111
`define OPC_Bcc		7'b1100011
`define OPC_Sx		7'b0100011

`endif

